* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 16 Feb 2013 05:47:49 PM CET

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

.temp 35.01

*Sheet Name:/
Lt 1 4 1.2uH
R1 1 3 12k
R2 3 0 3700
Cb 3 0 0.0033uF
Q1 4 3 6 Q2N3866
Re 6 7 44
LRFC 7 8 50uH
REE 8 0 700
CC 4 5 0.0033uF
C1 5 7 218pF
C2 7 0 2842pF IC=1V
Cf 5 0 20pF
RL 5 0 5371
ICC 1 0 -17
RICC 1 0 1
CICC 1 0 0.0033uF

.model Q2N3866 NPN (
+ IS = 9.798605E-15
+ BF = 145.568899
+ NF = 1.007933
+ VAF = 64.3030691
+ IKF = 0.3661244
+ ISE = 1.806705E-14
+ NE = 1.6207001
+ BR = 10.471
+ NR = 1.0003673
+ VAR = 8.322
+ IKR = 0.1449443
+ ISC = 3.326752E-15
+ NC = 1.1076801
+ RB = 15.986
+ IRB = 2.530217E-3
+ RBM = 0.01
+ RE = 0.02604
+ RC = 1.0359
+ CJE = 9.055532E-12
+ VJE = 0.6761546
+ MJE = 0.2754969
+ TF = 1.25476E-10
+ XTF = 13.0616413
+ VTF = 0.4699
+ ITF = 0.2828
+ PTF = 18.9645325
+ CJC = 7.054363E-12
+ VJC = 0.5769848
+ MJC = 0.3139067
+ XCJC = 1
+ TR = 5.698362E-8
+ CJS = 0
+ VJS = .75
+ MJS = 0
+ XTB = 1.831
+ EG = 1.11
+ XTI = 5.0205
+ KF = 0
+ AF = 1
+ FC = 0.9
+ )

.OP

.end

