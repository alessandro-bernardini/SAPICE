*low noise oscillator

ICC 0 1 12
RI 1 0 1
R1 1 2 10
Cbp1 2 0 0.2m
RCbp1 2 0 1000k
Q1 3 4 5 Q2N3866
LRFC1 5 6 100u
R2 6 0 47
Q2 8 7 5 Q2N3866
Ltrafo5 1 8 25u
Ltrafo6 10 0 25u
RLOAD 10 0 50
K1 Ltrafo5 Ltrafo6 0.99
Cbp2 7 0 0.1m
R3 7 0 1k
R4 1 7 3.9k
L1 2 3 0.05u
L3 4 7 0.05u
L2 9l 4 1.12u
RL2 9l 9 0.05
K2 L3 L2 0.99
K3 L1 L2 0.99
K4 L1 L3 0.99
C2 9 0 250p

.model Q2N3866 NPN (
+ IS = 9.798605E-15
+ BF = 145.568899
+ NF = 1.007933
+ VAF = 64.3030691
+ IKF = 0.3661244
+ ISE = 1.806705E-14
+ NE = 1.6207001
+ BR = 10.471
+ NR = 1.0003673
+ VAR = 8.322
+ IKR = 0.1449443
+ ISC = 3.326752E-15
+ NC = 1.1076801
+ RB = 15.986
+ IRB = 2.530217E-3
+ RBM = 0.01
+ RE = 0.02604
+ RC = 1.0359
+ CJE = 9.055532E-12
+ VJE = 0.6761546
+ MJE = 0.2754969
+ TF = 1.25476E-10
+ XTF = 13.0616413
+ VTF = 0.4699
+ ITF = 0.2828
+ PTF = 18.9645325
+ CJC = 7.054363E-12
+ VJC = 0.5769848
+ MJC = 0.3139067
+ XCJC = 1
+ TR = 5.698362E-8
+ CJS = 0
+ VJS = .75
+ MJS = 0
+ XTB = 1.831
+ EG = 1.11
+ XTI = 5.0205
+ KF = 0
+ AF = 1
+ FC = 0.9
+ )


