* simplest RLC example circuit

R1 1 0 1
L1 1 0 1H
C1 1 0 1
I1 1 0 1

.OP
.end
